** sch_path: /home/designer/shared/OS_AnalogIC_VLSISOC_Oct2025/design_data/transmission_gate.sch
**.subckt transmission_gate B GN GP A BP BN
*.iopin B
*.iopin GN
*.iopin A
*.iopin GP
*.iopin BN
*.iopin BP
XM1 A GN B BN sg13_lv_nmos w=10u l=0.13u ng=1 m=1
XM2 A GP B BP sg13_lv_pmos w=20u l=0.13u ng=2 m=1
**.ends
.end
